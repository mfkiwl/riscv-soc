//------------------------------------------------------------------------------
// Copyright 2022 Dominik Salvet
// https://github.com/dominiksalvet/riscv-soc
//------------------------------------------------------------------------------

module cpu (
    input rst_l,
    input clk
);
    
endmodule
